CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
177209362 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 587 600 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 45 526 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 138 268 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
12 Hex Display~
7 596 150 0 18 19
10 5 4 3 2 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6153 0 0
0
0
14 Logic Display~
6 1125 462 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
5 SCOPE
12 1074 476 0 1 11
0 2
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
14 Logic Display~
6 892 454 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
5 SCOPE
12 832 473 0 1 11
0 3
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 544 469 0 1 11
0 4
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
14 Logic Display~
6 596 456 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 288 454 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
12 SPDT Switch~
164 96 519 0 10 11
0 7 7 8 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8903 0 0
0
0
6 JK RN~
219 1028 506 0 6 22
0 10 3 10 6 11 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3834 0 0
0
0
6 JK RN~
219 742 503 0 6 22
0 10 4 10 6 12 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3363 0 0
0
0
6 JK RN~
219 466 498 0 6 22
0 10 5 10 6 13 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
7668 0 0
0
0
6 JK RN~
219 198 497 0 6 22
0 10 7 10 6 14 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
4718 0 0
0
0
5 SCOPE
12 246 467 0 1 11
0 5
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3874 0 0
0
0
5 SCOPE
12 125 471 0 1 11
0 7
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6671 0 0
0
0
7 Pulser~
4 64 418 0 10 12
0 15 16 7 17 0 0 5 5 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3789 0 0
0
0
32
0 4 2 0 0 8320 0 0 4 6 0 4
1059 489
1059 215
587 215
587 174
0 3 3 0 0 4224 0 0 4 9 0 4
791 486
791 204
593 204
593 174
0 2 4 0 0 4224 0 0 4 12 0 4
501 481
501 233
599 233
599 174
0 1 5 0 0 8320 0 0 4 14 0 4
228 480
228 189
605 189
605 174
1 0 2 0 0 0 0 6 0 0 6 2
1074 488
1074 489
6 1 2 0 0 0 0 13 5 0 0 3
1052 489
1125 489
1125 480
0 2 3 0 0 0 0 0 13 9 0 3
892 486
892 498
997 498
1 0 3 0 0 0 0 8 0 0 9 2
832 485
832 486
6 1 3 0 0 0 0 14 7 0 0 3
766 486
892 486
892 472
0 2 4 0 0 0 0 0 14 11 0 3
596 481
596 495
711 495
1 1 4 0 0 0 0 9 10 0 0 3
544 481
596 481
596 474
6 1 4 0 0 0 0 15 9 0 0 2
490 481
544 481
1 0 5 0 0 0 0 17 0 0 14 2
246 479
246 480
6 1 5 0 0 0 0 16 11 0 0 4
222 480
278 480
278 472
288 472
2 1 5 0 0 0 0 15 11 0 0 5
435 490
293 490
293 485
288 485
288 472
0 1 6 0 0 4096 0 0 1 19 0 2
588 553
588 587
4 0 6 0 0 0 0 15 0 0 19 2
466 529
466 553
4 0 6 0 0 0 0 14 0 0 19 2
742 534
742 553
4 4 6 0 0 8320 0 16 13 0 0 4
198 528
198 553
1028 553
1028 537
1 0 7 0 0 4096 0 18 0 0 21 2
125 483
125 489
1 2 7 0 0 8320 0 12 16 0 0 3
113 519
113 489
167 489
1 3 8 0 0 4224 0 2 12 0 0 4
57 526
71 526
71 523
79 523
3 2 7 0 0 8320 9 19 12 0 0 6
88 409
98 409
98 509
71 509
71 515
79 515
0 3 10 0 0 4096 0 0 16 25 0 3
168 480
168 498
174 498
0 1 10 0 0 4096 0 0 16 32 0 3
168 266
168 480
174 480
0 3 10 0 0 0 0 0 15 27 0 3
413 481
413 499
442 499
0 1 10 0 0 4096 0 0 15 32 0 3
413 266
413 481
442 481
0 3 10 0 0 0 0 0 14 30 0 3
705 486
705 504
718 504
1 0 10 0 0 0 0 3 0 0 32 2
150 268
150 268
0 1 10 0 0 4096 0 0 14 32 0 3
705 266
705 486
718 486
0 3 10 0 0 0 0 0 13 32 0 3
995 489
995 507
1004 507
0 1 10 0 0 8320 0 0 13 0 0 5
150 268
150 266
995 266
995 489
1004 489
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
