CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 303 448 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 160 451 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 186 329 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 866 330 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
5 SCOPE
12 830 322 0 1 11
0 4
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5394 0 0
0
0
9 2-In AND~
219 687 279 0 3 22
0 6 5 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7734 0 0
0
0
5 SCOPE
12 1044 320 0 1 11
0 7
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
14 Logic Display~
6 1086 313 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
6 JK RN~
219 987 350 0 6 22
0 3 10 3 9 13 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 3 0
1 U
3549 0 0
0
0
6 JK RN~
219 788 351 0 6 22
0 2 10 2 9 14 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 3 0
1 U
7931 0 0
0
0
5 SCOPE
12 141 333 0 1 11
0 10
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9325 0 0
0
0
12 SPDT Switch~
164 188 446 0 10 11
0 10 10 8 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8903 0 0
0
0
6 JK RN~
219 602 353 0 6 22
0 6 10 6 9 15 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
3834 0 0
0
0
5 SCOPE
12 499 325 0 1 11
0 6
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3363 0 0
0
0
9 2-In AND~
219 874 288 0 3 22
0 2 4 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -365013531
65 0 0 0 4 1 2 0
1 U
7668 0 0
0
0
14 Logic Display~
6 381 319 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
12 Hex Display~
7 596 176 0 18 19
10 6 5 4 7 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3874 0 0
0
0
7 Pulser~
4 130 392 0 10 12
0 16 17 10 18 0 0 5 5 4
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6671 0 0
0
0
6 JK RN~
219 314 353 0 6 22
0 12 10 12 9 19 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
3789 0 0
0
0
33
0 3 2 0 0 4096 0 0 10 2 0 3
753 334
753 352
764 352
0 1 2 0 0 4096 0 0 10 8 0 3
744 279
744 334
764 334
1 3 3 0 0 8192 0 9 9 0 0 4
963 333
953 333
953 351
963 351
3 1 3 0 0 4224 0 15 9 0 0 3
895 288
963 288
963 333
1 0 4 0 0 0 0 4 0 0 7 2
850 334
850 334
1 0 4 0 0 0 0 5 0 0 7 2
830 334
830 334
6 2 4 0 0 4096 0 10 15 0 0 3
812 334
850 334
850 297
3 1 2 0 0 4224 0 6 15 0 0 2
708 279
850 279
0 2 5 0 0 8192 0 0 6 13 0 3
626 287
626 288
663 288
0 1 6 0 0 8192 0 0 6 31 0 3
535 336
535 270
663 270
1 0 7 0 0 4096 0 7 0 0 12 2
1044 332
1044 331
6 1 7 0 0 8192 0 9 8 0 0 3
1011 333
1011 331
1086 331
6 2 5 0 0 4224 0 13 17 0 0 4
626 336
626 264
599 264
599 200
6 3 4 0 0 8320 0 10 17 0 0 4
812 334
812 239
593 239
593 200
6 4 7 0 0 8320 0 9 17 0 0 4
1011 333
1011 214
587 214
587 200
1 3 8 0 0 4224 0 2 12 0 0 3
172 451
172 450
171 450
1 0 9 0 0 4096 0 1 0 0 20 2
315 448
314 448
0 4 9 0 0 4096 0 0 13 20 0 4
603 449
603 392
602 392
602 384
0 4 9 0 0 4096 0 0 10 20 0 2
788 449
788 382
4 4 9 0 0 8320 0 19 9 0 0 4
314 384
314 449
987 449
987 381
0 2 10 0 0 4096 0 0 13 23 0 3
521 420
521 345
571 345
0 2 10 0 0 4096 0 0 10 23 0 3
718 420
718 343
757 343
0 2 10 0 0 4224 0 0 9 25 0 4
205 420
942 420
942 342
956 342
0 1 10 0 0 0 0 0 11 25 0 2
205 345
141 345
1 2 10 0 0 0 0 12 19 0 0 3
205 446
205 345
283 345
3 2 10 0 0 8320 11 18 12 0 0 4
154 383
165 383
165 442
171 442
0 3 6 0 0 0 0 0 13 31 0 3
557 336
557 354
578 354
0 1 6 0 0 8192 0 0 17 31 0 4
436 336
436 208
605 208
605 200
1 0 6 0 0 0 0 16 0 0 31 2
381 337
381 336
1 0 6 0 0 0 0 14 0 0 31 2
499 337
499 336
6 1 6 0 0 4224 0 19 13 0 0 2
338 336
578 336
0 3 12 0 0 4096 0 0 19 33 0 3
275 336
275 354
290 354
1 1 12 0 0 4224 0 3 19 0 0 4
198 329
275 329
275 336
290 336
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
