CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 617 566 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 167 691 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 45 526 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 138 268 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
9 2-In AND~
219 888 588 0 3 22
0 6 7 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 6 0
1 U
5394 0 0
0
0
8 2-In OR~
219 957 618 0 3 22
0 9 8 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 4 0
1 U
7734 0 0
0
0
9 2-In AND~
219 885 649 0 3 22
0 2 5 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
9914 0 0
0
0
9 Inverter~
13 839 619 0 2 22
0 2 7
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 5 0
1 U
3747 0 0
0
0
9 2-In AND~
219 600 597 0 3 22
0 11 12 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
3549 0 0
0
0
8 2-In OR~
219 672 636 0 3 22
0 14 13 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 4 0
1 U
7931 0 0
0
0
9 2-In AND~
219 600 666 0 3 22
0 2 10 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
9325 0 0
0
0
9 Inverter~
13 552 628 0 2 22
0 2 12
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 5 0
1 U
8903 0 0
0
0
9 2-In AND~
219 318 583 0 3 22
0 17 19 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
3834 0 0
0
0
8 2-In OR~
219 387 613 0 3 22
0 21 20 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 4 0
1 U
3363 0 0
0
0
9 2-In AND~
219 315 644 0 3 22
0 2 16 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
7668 0 0
0
0
9 Inverter~
13 269 614 0 2 22
0 2 19
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 5 0
1 U
4718 0 0
0
0
12 Hex Display~
7 596 150 0 18 19
10 17 11 6 22 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3874 0 0
0
0
14 Logic Display~
6 1125 462 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
5 SCOPE
12 1074 476 0 1 11
0 22
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3789 0 0
0
0
14 Logic Display~
6 892 454 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
5 SCOPE
12 832 473 0 1 11
0 6
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3750 0 0
0
0
5 SCOPE
12 544 469 0 1 11
0 11
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8778 0 0
0
0
14 Logic Display~
6 596 456 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 288 454 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
12 SPDT Switch~
164 96 519 0 10 11
0 23 23 24 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3136 0 0
0
0
6 JK RN~
219 1028 506 0 6 22
0 26 4 26 15 27 22
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
5950 0 0
0
0
6 JK RN~
219 742 503 0 6 22
0 26 3 26 15 5 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
5670 0 0
0
0
6 JK RN~
219 466 498 0 6 22
0 26 18 26 15 10 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
6828 0 0
0
0
6 JK RN~
219 198 497 0 6 22
0 26 23 26 15 16 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
6735 0 0
0
0
5 SCOPE
12 246 467 0 1 11
0 17
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8365 0 0
0
0
5 SCOPE
12 125 471 0 1 11
0 23
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4132 0 0
0
0
7 Pulser~
4 64 418 0 10 12
0 28 29 23 30 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4551 0 0
0
0
53
0 0 2 0 0 4096 0 0 0 3 22 2
272 692
272 635
0 0 2 0 0 0 0 0 0 3 14 4
557 692
557 678
555 678
555 656
1 0 2 0 0 8336 0 2 0 0 8 4
179 691
179 692
852 692
852 640
3 2 3 0 0 8320 0 10 27 0 0 3
705 636
711 636
711 495
3 2 4 0 0 8320 0 6 26 0 0 3
990 618
997 618
997 498
2 5 5 0 0 8320 0 7 27 0 0 4
861 658
798 658
798 504
772 504
1 0 6 0 0 8192 0 5 0 0 33 3
864 579
808 579
808 486
1 1 2 0 0 0 0 8 7 0 0 3
842 637
842 640
861 640
2 2 7 0 0 8320 0 8 5 0 0 3
842 601
842 597
864 597
3 2 8 0 0 4224 0 7 6 0 0 4
906 649
936 649
936 627
944 627
3 1 9 0 0 4224 0 5 6 0 0 4
909 588
936 588
936 609
944 609
2 5 10 0 0 8320 0 11 28 0 0 4
576 675
511 675
511 499
496 499
1 0 11 0 0 8192 0 9 0 0 35 3
576 588
521 588
521 481
1 1 2 0 0 0 0 12 11 0 0 3
555 646
555 657
576 657
2 2 12 0 0 8320 0 12 9 0 0 3
555 610
555 606
576 606
3 2 13 0 0 4224 0 11 10 0 0 4
621 666
649 666
649 645
659 645
3 1 14 0 0 8320 0 9 10 0 0 4
621 597
649 597
649 627
659 627
1 0 15 0 0 0 0 1 0 0 40 2
618 553
618 553
2 5 16 0 0 8320 0 15 29 0 0 3
291 653
228 653
228 498
1 0 17 0 0 8192 0 13 0 0 37 3
294 574
238 574
238 480
3 2 18 0 0 4224 0 14 28 0 0 3
420 613
420 490
435 490
1 1 2 0 0 0 0 16 15 0 0 3
272 632
272 635
291 635
2 2 19 0 0 8320 0 16 13 0 0 3
272 596
272 592
294 592
3 2 20 0 0 4224 0 15 14 0 0 4
336 644
366 644
366 622
374 622
3 1 21 0 0 4224 0 13 14 0 0 4
339 583
366 583
366 604
374 604
0 4 22 0 0 8320 0 0 17 31 0 4
1059 489
1059 215
587 215
587 174
0 3 6 0 0 4224 0 0 17 33 0 4
791 486
791 204
593 204
593 174
0 2 11 0 0 4224 0 0 17 35 0 4
501 481
501 233
599 233
599 174
0 1 17 0 0 8320 0 0 17 37 0 4
228 480
228 189
605 189
605 174
1 0 22 0 0 0 0 19 0 0 31 2
1074 488
1074 489
6 1 22 0 0 0 0 26 18 0 0 3
1052 489
1125 489
1125 480
1 0 6 0 0 0 0 21 0 0 33 2
832 485
832 486
6 1 6 0 0 0 0 27 20 0 0 3
766 486
892 486
892 472
1 1 11 0 0 0 0 22 23 0 0 3
544 481
596 481
596 474
6 1 11 0 0 0 0 28 22 0 0 2
490 481
544 481
1 0 17 0 0 0 0 30 0 0 37 2
246 479
246 480
6 1 17 0 0 0 0 29 24 0 0 4
222 480
278 480
278 472
288 472
4 0 15 0 0 4096 0 28 0 0 40 2
466 529
466 553
4 0 15 0 0 0 0 27 0 0 40 2
742 534
742 553
4 4 15 0 0 8320 0 29 26 0 0 4
198 528
198 553
1028 553
1028 537
1 0 23 0 0 4096 0 31 0 0 42 2
125 483
125 489
1 2 23 0 0 8320 0 25 29 0 0 3
113 519
113 489
167 489
1 3 24 0 0 4224 0 3 25 0 0 4
57 526
71 526
71 523
79 523
3 2 23 0 0 8320 25 32 25 0 0 6
88 409
98 409
98 509
71 509
71 515
79 515
0 3 26 0 0 4096 0 0 29 46 0 3
168 480
168 498
174 498
0 1 26 0 0 4096 0 0 29 53 0 3
168 266
168 480
174 480
0 3 26 0 0 0 0 0 28 48 0 3
413 481
413 499
442 499
0 1 26 0 0 4096 0 0 28 53 0 3
413 266
413 481
442 481
0 3 26 0 0 0 0 0 27 51 0 3
705 486
705 504
718 504
1 0 26 0 0 0 0 4 0 0 53 2
150 268
150 268
0 1 26 0 0 4096 0 0 27 53 0 3
705 266
705 486
718 486
0 3 26 0 0 0 0 0 26 53 0 3
995 489
995 507
1004 507
0 1 26 0 0 8320 0 0 26 0 0 5
150 268
150 266
995 266
995 489
1004 489
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
