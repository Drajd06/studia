CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 16 523 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 617 566 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 138 268 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
5 SCOPE
12 1250 179 0 1 11
0 4
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
10 2-In NAND~
219 1147 192 0 3 22
0 2 3 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1703441668
65 0 0 0 4 1 3 0
1 U
5394 0 0
0
0
9 2-In AND~
219 138 488 0 3 22
0 5 4 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2122937626
65 0 0 0 4 1 4 0
1 U
7734 0 0
0
0
7 Pulser~
4 35 415 0 10 12
0 13 14 5 15 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9914 0 0
0
0
5 SCOPE
12 95 467 0 1 11
0 5
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
12 SPDT Switch~
164 67 516 0 10 11
0 5 5 7 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3549 0 0
0
0
12 Hex Display~
7 596 150 0 18 19
10 2 9 3 11 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7931 0 0
0
0
14 Logic Display~
6 1125 462 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
5 SCOPE
12 1074 476 0 1 11
0 11
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8903 0 0
0
0
14 Logic Display~
6 892 454 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
5 SCOPE
12 832 473 0 1 11
0 3
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 544 469 0 1 11
0 9
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7668 0 0
0
0
14 Logic Display~
6 596 456 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 288 454 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
6 JK RN~
219 1028 506 0 6 22
0 12 3 12 10 16 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
6671 0 0
0
0
6 JK RN~
219 742 503 0 6 22
0 12 9 12 10 17 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3789 0 0
0
0
6 JK RN~
219 466 498 0 6 22
0 12 2 12 10 18 9
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
4871 0 0
0
0
6 JK RN~
219 198 497 0 6 22
0 12 6 12 10 19 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
3750 0 0
0
0
5 SCOPE
12 246 467 0 1 11
0 2
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8778 0 0
0
0
37
0 1 2 0 0 8320 0 0 5 12 0 5
344 490
344 96
1103 96
1103 183
1123 183
0 2 3 0 0 4224 0 0 5 5 0 3
949 498
949 201
1123 201
0 1 4 0 0 8192 0 0 4 4 0 3
1218 193
1218 191
1250 191
2 3 4 0 0 8320 0 6 5 0 0 5
114 497
114 625
1218 625
1218 192
1174 192
0 2 3 0 0 0 0 0 18 21 0 3
892 486
892 498
997 498
1 0 5 0 0 0 0 8 0 0 7 2
95 479
95 479
1 1 5 0 0 4224 0 9 6 0 0 3
84 516
84 479
114 479
3 2 6 0 0 8320 0 6 21 0 0 3
159 488
159 489
167 489
1 3 7 0 0 4224 0 1 9 0 0 4
28 523
42 523
42 520
50 520
3 2 5 0 0 8320 8 7 9 0 0 6
59 406
69 406
69 506
42 506
42 512
50 512
0 2 9 0 0 8192 0 0 19 22 0 3
595 481
595 495
711 495
1 2 2 0 0 0 0 17 20 0 0 3
288 472
288 490
435 490
1 0 10 0 0 0 0 2 0 0 28 2
618 553
618 553
0 4 11 0 0 8320 0 0 10 19 0 4
1059 489
1059 215
587 215
587 174
0 3 3 0 0 128 0 0 10 21 0 4
791 486
791 204
593 204
593 174
0 2 9 0 0 4224 0 0 10 23 0 4
501 481
501 233
599 233
599 174
0 1 2 0 0 128 0 0 10 25 0 4
228 480
228 189
605 189
605 174
1 0 11 0 0 0 0 12 0 0 19 2
1074 488
1074 489
6 1 11 0 0 0 0 18 11 0 0 3
1052 489
1125 489
1125 480
1 0 3 0 0 0 0 14 0 0 21 2
832 485
832 486
6 1 3 0 0 0 0 19 13 0 0 3
766 486
892 486
892 472
1 1 9 0 0 0 0 15 16 0 0 3
544 481
596 481
596 474
6 1 9 0 0 0 0 20 15 0 0 2
490 481
544 481
1 0 2 0 0 0 0 22 0 0 25 2
246 479
246 480
6 1 2 0 0 0 0 21 17 0 0 4
222 480
278 480
278 472
288 472
4 0 10 0 0 4096 0 20 0 0 28 2
466 529
466 553
4 0 10 0 0 0 0 19 0 0 28 2
742 534
742 553
4 4 10 0 0 8320 0 21 18 0 0 4
198 528
198 553
1028 553
1028 537
0 3 12 0 0 4096 0 0 21 30 0 3
168 480
168 498
174 498
0 1 12 0 0 4096 0 0 21 37 0 3
168 266
168 480
174 480
0 3 12 0 0 0 0 0 20 32 0 3
413 481
413 499
442 499
0 1 12 0 0 4096 0 0 20 37 0 3
413 266
413 481
442 481
0 3 12 0 0 0 0 0 19 35 0 3
705 486
705 504
718 504
1 0 12 0 0 0 0 3 0 0 37 2
150 268
150 268
0 1 12 0 0 4096 0 0 19 37 0 3
705 266
705 486
718 486
0 3 12 0 0 0 0 0 18 37 0 3
995 489
995 507
1004 507
0 1 12 0 0 8320 0 0 18 0 0 5
150 268
150 266
995 266
995 489
1004 489
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
