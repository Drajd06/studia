CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 645 1872 1004
193986578 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 691 411 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V17
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 509 300 0 1 11
0 16
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V16
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 689 576 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V15
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 508 429 0 1 11
0 5
0
0 0 21360 90
2 0V
11 0 25 8
3 V14
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 277 402 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V13
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 255 656 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 210 303 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 830 78 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 829 214 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 765 119 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 597 104 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 596 222 0 1 11
0 25
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 525 135 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 341 194 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 257 75 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 260 160 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4718 0 0
0
0
5 SCOPE
12 375 449 0 1 11
0 3
0
0 0 57584 0
3 TP9
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3874 0 0
0
0
5 SCOPE
12 442 550 0 1 11
0 2
0
0 0 57584 0
3 TP7
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6671 0 0
0
0
5 SCOPE
12 775 439 0 1 11
0 12
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3789 0 0
0
0
5 SCOPE
12 602 331 0 1 11
0 13
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4871 0 0
0
0
5 SCOPE
12 330 294 0 1 11
0 14
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3750 0 0
0
0
14 Logic Display~
6 396 539 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 411 425 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 830 431 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 648 320 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 362 286 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5950 0 0
0
0
6 JK RN~
219 257 589 0 6 22
0 7 4 2 6 7 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 6 0
1 U
5670 0 0
0
0
12 D Flip-Flop~
219 307 514 0 4 9
0 11 4 11 3
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
6828 0 0
0
0
5 7474~
219 691 506 0 6 22
0 10 8 4 15 8 12
0
0 0 4720 0
6 74LS74
0 -60 42 -52
3 U6A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 0 2 1 5 0
1 U
6735 0 0
0
0
5 4013~
219 509 396 0 6 22
0 16 9 4 5 9 13
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 0 2 1 4 0
1 U
8365 0 0
0
0
6 JK RN~
219 278 334 0 6 22
0 18 4 18 17 31 14
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
4132 0 0
0
0
5 SCOPE
12 901 105 0 1 11
0 19
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4551 0 0
0
0
14 Logic Display~
6 945 85 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3635 0 0
0
0
5 SCOPE
12 657 126 0 1 11
0 23
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3973 0 0
0
0
14 Logic Display~
6 694 114 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3851 0 0
0
0
14 Logic Display~
6 435 72 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8383 0 0
0
0
6 74112~
219 830 169 0 7 32
0 21 22 4 22 20 32 19
0
0 0 4720 0
7 74LS112
-3 -60 46 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 467298223
65 0 0 512 2 1 3 0
1 U
9334 0 0
0
0
5 4027~
219 597 191 0 7 32
0 24 26 4 26 25 33 23
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 215639992
65 0 0 512 2 1 2 0
1 U
7471 0 0
0
0
6 JK RN~
219 342 132 0 6 22
0 29 4 28 27 34 30
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
3334 0 0
0
0
5 SCOPE
12 398 92 0 1 11
0 30
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3559 0 0
0
0
5 SCOPE
12 222 93 0 1 11
0 4
0
0 0 57584 0
3 TP8
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
984 0 0
0
0
7 Pulser~
4 130 133 0 10 12
0 35 36 4 37 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7557 0 0
0
0
49
0 1 2 0 0 4096 0 0 18 6 0 3
396 572
442 572
442 562
0 1 3 0 0 4096 0 0 17 16 0 4
376 478
376 469
375 469
375 461
1 0 4 0 0 4096 0 41 0 0 47 2
222 105
222 124
1 4 5 0 0 4224 0 4 30 0 0 2
509 416
509 402
6 0 2 0 0 4096 0 27 0 0 6 2
281 572
354 572
3 1 2 0 0 8320 0 27 22 0 0 6
233 590
233 630
354 630
354 572
396 572
396 557
1 4 6 0 0 4224 0 6 27 0 0 4
256 643
256 628
257 628
257 620
1 5 7 0 0 8320 0 27 27 0 0 5
233 572
233 536
308 536
308 590
287 590
2 5 8 0 0 8320 0 29 29 0 0 5
667 470
667 436
730 436
730 488
721 488
2 5 9 0 0 8320 0 30 30 0 0 5
485 360
485 328
548 328
548 378
539 378
0 3 4 0 0 8192 0 0 29 13 0 3
468 378
468 488
667 488
1 1 10 0 0 4224 0 29 1 0 0 2
691 443
691 423
0 3 4 0 0 0 0 0 30 43 0 4
166 431
352 431
352 378
485 378
0 2 4 0 0 0 0 0 28 43 0 2
166 496
283 496
1 3 11 0 0 8320 0 28 28 0 0 5
283 478
283 452
351 452
351 496
337 496
4 1 3 0 0 4224 0 28 23 0 0 3
331 478
411 478
411 443
0 1 12 0 0 4096 0 0 19 19 0 2
775 470
775 451
0 1 13 0 0 4096 0 0 20 20 0 2
602 360
602 343
6 1 12 0 0 4224 0 29 24 0 0 3
715 470
830 470
830 449
6 1 13 0 0 4224 0 30 25 0 0 3
533 360
648 360
648 338
0 1 14 0 0 12288 0 0 21 22 0 4
331 317
331 314
330 314
330 306
6 1 14 0 0 4224 0 31 26 0 0 3
302 317
362 317
362 304
4 1 15 0 0 4224 0 29 3 0 0 4
691 518
691 548
690 548
690 563
1 1 16 0 0 4224 0 2 30 0 0 2
509 312
509 339
4 1 17 0 0 4224 0 31 5 0 0 2
278 365
278 389
0 3 18 0 0 4224 0 0 31 28 0 3
239 315
239 335
254 335
0 2 4 0 0 0 0 0 31 43 0 2
166 326
247 326
1 1 18 0 0 0 0 7 31 0 0 4
222 303
239 303
239 317
254 317
1 0 19 0 0 4096 0 32 0 0 30 2
901 117
901 133
7 1 19 0 0 4224 0 37 33 0 0 3
854 133
945 133
945 103
1 5 20 0 0 4224 0 9 37 0 0 2
830 201
830 181
1 1 21 0 0 4224 0 37 8 0 0 2
830 106
830 90
0 4 22 0 0 4224 0 0 37 34 0 3
800 133
800 151
806 151
1 2 22 0 0 0 0 10 37 0 0 4
777 119
792 119
792 133
806 133
0 3 4 0 0 4096 0 0 37 42 0 4
546 250
781 250
781 142
800 142
0 1 23 0 0 4096 0 0 34 37 0 2
657 155
657 138
7 1 23 0 0 4224 0 38 35 0 0 3
621 155
694 155
694 132
1 1 24 0 0 4224 0 11 38 0 0 2
597 116
597 134
1 5 25 0 0 4224 0 12 38 0 0 2
597 209
597 197
0 4 26 0 0 4096 0 0 38 41 0 3
565 155
565 173
573 173
1 2 26 0 0 4224 0 13 38 0 0 4
537 135
565 135
565 155
573 155
0 3 4 0 0 4096 0 0 38 43 0 4
166 250
546 250
546 164
573 164
0 2 4 0 0 4224 0 0 27 47 0 3
166 124
166 581
226 581
1 4 27 0 0 4224 0 14 39 0 0 2
342 181
342 163
1 3 28 0 0 4224 0 16 39 0 0 4
272 160
303 160
303 133
318 133
1 1 29 0 0 8320 0 15 39 0 0 4
269 75
303 75
303 115
318 115
3 2 4 0 0 0 0 42 39 0 0 2
154 124
311 124
0 1 30 0 0 4096 0 0 40 49 0 2
398 115
398 104
6 1 30 0 0 4224 0 39 36 0 0 3
366 115
435 115
435 90
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
243 428 339 449
251 435 339 450
11 narastajace
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
240 258 320 279
248 264 320 279
9 opadajaca
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
714 394 810 415
722 401 810 416
11 narastajace
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
529 287 625 308
537 294 625 309
11 narastajace
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
224 512 304 533
232 518 304 533
9 opadajaca
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
788 17 868 38
796 23 868 38
9 opadajaca
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
545 45 641 66
553 52 641 67
11 narastajace
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
308 50 388 71
316 56 388 71
9 opadajaca
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
