CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 1 120 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 1040
143654930 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 375 215 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 301 474 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 160 451 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 186 329 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
12 D Flip-Flop~
219 1153 214 0 4 9
0 2 2 23 3
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U12
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
9 2-In AND~
219 995 98 0 3 22
0 5 4 2
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U11A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 7 0
1 U
7734 0 0
0
0
14 Logic Display~
6 1074 301 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
6 JK RN~
219 1015 335 0 6 22
0 13 7 13 9 24 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 U10A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 6 0
1 U
3747 0 0
0
0
8 2-In OR~
219 900 327 0 3 22
0 15 14 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
9 3-In AND~
219 837 367 0 4 22
0 8 6 3 14
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 5 0
1 U
7931 0 0
0
0
9 3-In AND~
219 839 296 0 4 22
0 10 5 11 15
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
9325 0 0
0
0
9 Inverter~
13 425 201 0 2 22
0 3 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
8903 0 0
0
0
5 SCOPE
12 498 108 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 449 108 0 1 11
0 11
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 380 112 0 1 11
0 5
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
12 Hex Display~
7 292 88 0 18 19
10 5 11 4 12 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4718 0 0
0
0
6 JK RN~
219 718 346 0 6 22
0 16 7 16 9 8 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
3874 0 0
0
0
8 2-In OR~
219 563 338 0 3 22
0 18 17 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -516008466
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
9 2-In AND~
219 487 372 0 3 22
0 6 3 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
3789 0 0
0
0
9 2-In AND~
219 486 312 0 3 22
0 10 5 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
4871 0 0
0
0
5 SCOPE
12 141 333 0 1 11
0 7
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
12 SPDT Switch~
164 188 446 0 10 11
0 7 7 19 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8778 0 0
0
0
14 Logic Display~
6 364 318 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
7 Pulser~
4 130 392 0 10 12
0 25 26 7 27 0 0 5 5 2
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6843 0 0
0
0
6 JK RN~
219 314 353 0 6 22
0 21 7 21 9 6 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3136 0 0
0
0
45
3 1 2 0 0 4224 0 6 5 0 0 3
994 74
1129 74
1129 178
3 2 4 0 0 4096 0 0 6 27 0 2
1003 135
1003 119
1 1 5 0 0 4096 0 0 6 27 0 2
985 135
985 119
0 2 6 0 0 8320 0 0 10 37 0 5
428 354
428 394
797 394
797 367
813 367
0 2 7 0 0 4096 0 0 8 32 0 3
686 428
984 428
984 327
0 2 3 0 0 0 0 0 19 7 0 2
463 414
463 381
1 3 3 0 0 128 0 12 10 0 0 4
410 201
410 414
813 414
813 376
5 1 8 0 0 4224 0 17 10 0 0 3
748 347
813 347
813 358
1 0 9 0 0 4096 0 2 0 0 11 2
313 474
314 473
0 4 9 0 0 8192 0 0 17 11 0 3
719 473
718 473
718 377
4 4 9 0 0 8320 0 25 8 0 0 4
314 384
314 473
1015 473
1015 366
0 2 5 0 0 8320 0 0 11 36 0 3
428 336
428 296
815 296
0 1 10 0 0 4096 0 0 20 15 0 3
458 201
458 303
462 303
0 3 11 0 0 4096 0 0 11 17 0 3
763 329
815 329
815 305
2 1 10 0 0 4224 0 12 11 0 0 3
446 201
815 201
815 287
0 1 5 0 0 0 0 0 0 36 27 2
347 336
347 135
6 2 11 0 0 8320 0 17 0 0 27 3
742 329
763 329
763 135
0 1 4 0 0 8192 0 0 7 19 0 3
1050 318
1050 319
1074 319
6 3 4 0 0 8320 0 8 0 0 27 3
1039 318
1050 318
1050 135
3 1 4 0 0 0 0 0 13 27 0 4
499 135
499 128
498 128
498 120
2 1 11 0 0 0 0 0 14 27 0 2
449 135
449 120
1 1 5 0 0 0 0 0 15 27 0 2
380 135
380 124
4 4 12 0 0 4224 0 0 16 27 0 2
283 135
283 112
3 3 4 0 0 0 0 0 16 27 0 2
289 135
289 112
2 2 11 0 0 0 0 0 16 27 0 2
295 135
295 112
1 1 5 0 0 0 0 0 16 27 0 2
301 135
301 112
-6369869 0 1 0 0 4256 0 0 0 0 0 2
250 135
1058 135
0 3 13 0 0 8192 0 0 8 29 0 3
969 327
969 336
991 336
3 1 13 0 0 4224 0 9 8 0 0 4
933 327
969 327
969 318
991 318
4 2 14 0 0 8320 0 10 9 0 0 4
858 367
879 367
879 336
887 336
4 1 15 0 0 8320 0 11 9 0 0 4
860 296
879 296
879 318
887 318
0 2 7 0 0 4224 0 0 17 42 0 3
205 428
687 428
687 338
0 3 16 0 0 8192 0 0 17 34 0 3
678 338
678 347
694 347
3 1 16 0 0 4224 0 18 17 0 0 4
596 338
678 338
678 329
694 329
1 0 5 0 0 0 0 23 0 0 36 2
364 336
364 336
6 2 5 0 0 0 0 25 20 0 0 4
338 336
455 336
455 321
462 321
5 1 6 0 0 0 0 25 19 0 0 4
344 354
455 354
455 363
463 363
3 2 17 0 0 4224 0 19 18 0 0 3
508 372
550 372
550 347
3 1 18 0 0 4224 0 20 18 0 0 3
507 312
550 312
550 329
1 3 19 0 0 4224 0 3 22 0 0 3
172 451
172 450
171 450
0 1 7 0 0 0 0 0 21 42 0 2
205 345
141 345
1 2 7 0 0 0 0 22 25 0 0 3
205 446
205 345
283 345
3 2 7 0 0 8320 20 24 22 0 0 4
154 383
165 383
165 442
171 442
0 3 21 0 0 4096 0 0 25 45 0 3
275 336
275 354
290 354
1 1 21 0 0 4224 0 4 25 0 0 4
198 329
275 329
275 336
290 336
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
