CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 1 120 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 1004
143654930 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 589 643 0 1 11
0 4
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 617 566 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 45 526 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 138 268 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
9 2-In XOR~
219 646 493 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 950 493 0 3 22
0 6 4 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 336 491 0 3 22
0 7 4 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -2122938140
65 0 0 0 4 1 3 0
1 U
9914 0 0
0
0
12 Hex Display~
7 596 150 0 18 19
10 7 5 6 10 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3747 0 0
0
0
14 Logic Display~
6 1125 462 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
5 SCOPE
12 1074 476 0 1 11
0 10
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
14 Logic Display~
6 892 454 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
5 SCOPE
12 832 473 0 1 11
0 6
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 544 469 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3834 0 0
0
0
14 Logic Display~
6 596 456 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 288 454 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
12 SPDT Switch~
164 96 519 0 10 11
0 11 11 12 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
4718 0 0
0
0
6 JK RN~
219 1028 506 0 6 22
0 14 2 14 9 16 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3874 0 0
0
0
6 JK RN~
219 742 503 0 6 22
0 14 3 14 9 17 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
6671 0 0
0
0
6 JK RN~
219 466 498 0 6 22
0 14 8 14 9 18 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
3789 0 0
0
0
6 JK RN~
219 198 497 0 6 22
0 14 11 14 9 19 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
4871 0 0
0
0
5 SCOPE
12 246 467 0 1 11
0 7
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3750 0 0
0
0
5 SCOPE
12 125 471 0 1 11
0 11
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8778 0 0
0
0
7 Pulser~
4 64 418 0 10 12
0 20 21 11 22 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
538 0 0
0
0
38
3 2 2 0 0 12416 0 6 17 0 0 4
983 493
989 493
989 498
997 498
3 2 3 0 0 4224 0 5 18 0 0 4
679 493
703 493
703 495
711 495
1 0 4 0 0 4096 0 1 0 0 5 2
590 630
591 630
1 0 5 0 0 4096 0 5 0 0 19 3
630 484
596 484
596 481
0 2 4 0 0 4096 0 0 5 7 0 3
591 630
591 502
630 502
1 0 6 0 0 4096 0 6 0 0 18 3
934 484
892 484
892 486
2 2 4 0 0 8320 0 7 6 0 0 5
320 500
320 630
923 630
923 502
934 502
1 1 7 0 0 8192 0 15 7 0 0 3
288 472
288 482
320 482
3 2 8 0 0 4224 0 7 19 0 0 4
369 491
427 491
427 490
435 490
1 0 9 0 0 0 0 2 0 0 25 2
618 553
618 553
0 4 10 0 0 8320 0 0 8 16 0 4
1059 489
1059 215
587 215
587 174
0 3 6 0 0 4224 0 0 8 18 0 4
791 486
791 204
593 204
593 174
0 2 5 0 0 4224 0 0 8 20 0 4
501 481
501 233
599 233
599 174
0 1 7 0 0 8320 0 0 8 22 0 4
228 480
228 189
605 189
605 174
1 0 10 0 0 0 0 10 0 0 16 2
1074 488
1074 489
6 1 10 0 0 0 0 17 9 0 0 3
1052 489
1125 489
1125 480
1 0 6 0 0 0 0 12 0 0 18 2
832 485
832 486
6 1 6 0 0 0 0 18 11 0 0 3
766 486
892 486
892 472
1 1 5 0 0 0 0 13 14 0 0 3
544 481
596 481
596 474
6 1 5 0 0 0 0 19 13 0 0 2
490 481
544 481
1 0 7 0 0 0 0 21 0 0 22 2
246 479
246 480
6 1 7 0 0 0 0 20 15 0 0 4
222 480
278 480
278 472
288 472
4 0 9 0 0 4096 0 19 0 0 25 2
466 529
466 553
4 0 9 0 0 0 0 18 0 0 25 2
742 534
742 553
4 4 9 0 0 8320 0 20 17 0 0 4
198 528
198 553
1028 553
1028 537
1 0 11 0 0 4096 0 22 0 0 27 2
125 483
125 489
1 2 11 0 0 8320 0 16 20 0 0 3
113 519
113 489
167 489
1 3 12 0 0 4224 0 3 16 0 0 4
57 526
71 526
71 523
79 523
3 2 11 0 0 8320 13 23 16 0 0 6
88 409
98 409
98 509
71 509
71 515
79 515
0 3 14 0 0 4096 0 0 20 31 0 3
168 480
168 498
174 498
0 1 14 0 0 4096 0 0 20 38 0 3
168 266
168 480
174 480
0 3 14 0 0 0 0 0 19 33 0 3
413 481
413 499
442 499
0 1 14 0 0 4096 0 0 19 38 0 3
413 266
413 481
442 481
0 3 14 0 0 0 0 0 18 36 0 3
705 486
705 504
718 504
1 0 14 0 0 0 0 4 0 0 38 2
150 268
150 268
0 1 14 0 0 4096 0 0 18 38 0 3
705 266
705 486
718 486
0 3 14 0 0 0 0 0 17 38 0 3
995 489
995 507
1004 507
0 1 14 0 0 8320 0 0 17 0 0 5
150 268
150 266
995 266
995 489
1004 489
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
